module PRNO_tb;
  reg clk_tb;
  reg [0:9] ao, bo;
  wire [0:1799] po;
  wire [0:23] fo, lo;
reg  [0:9]r0[0:64];
reg [0:9]r1[0:64];
integer i;

  PRNO P(.clk(clk_tb), .R0_in(ao), .R1_in(bo), .P(po), .first(fo), .last(lo));

initial
begin
    clk_tb = 0;
end

always
begin
    #5;
    clk_tb = ~ clk_tb;
end


  initial begin
r0[0 ]=10'b0110111011;
r0[1 ]=10'b0111101000;
r0[2 ]=10'b1100000001;
r0[3 ]=10'b0110110110;
r0[4 ]=10'b0100011000;
r0[5 ]=10'b0011111100;
r0[6 ]=10'b0011111100;
r0[7 ]=10'b1111000101;
r0[8 ]=10'b0011001100;
r0[9 ]=10'b1000011010;
r0[10]=10'b0001001001;
r0[11]=10'b0110101011;
r0[12]=10'b0101110000;
r0[13]=10'b0010110011;
r0[14]=10'b1110000111;
r0[15]=10'b1000000000;
r0[16]=10'b1111101101;
r0[17]=10'b1111101011;
r0[18]=10'b0010001011;
r0[19]=10'b0011101000;
r0[20]=10'b0011011010;
r0[21]=10'b0011111100;
r0[22]=10'b0111001100;
r0[23]=10'b1000101110;
r0[24]=10'b0101000010;
r0[25]=10'b0000101010;
r0[26]=10'b0000100001;
r0[27]=10'b1000010000;
r0[28]=10'b1011100100;
r0[29]=10'b0110111111;
r0[30]=10'b1001110000;
r0[31]=10'b1101110101;
r0[32]=10'b0101111100;
r0[33]=10'b1011001000;
r0[34]=10'b1000001100;
r0[35]=10'b0001100101;
r0[36]=10'b0000000010;
r0[37]=10'b0010100011;
r0[38]=10'b1111010010;
r0[39]=10'b0000100101;
r0[40]=10'b0100111011;
r0[41]=10'b0110111001;
r0[42]=10'b0010011101;
r0[43]=10'b1000011010;
r0[44]=10'b0010000010;
r0[45]=10'b1001001111;
r0[46]=10'b1111001111;
r0[47]=10'b0010110010;
r0[48]=10'b0111111110;
r0[49]=10'b0100100011;
r0[50]=10'b0100001110;
r0[51]=10'b0111101101;
r0[52]=10'b1000010010;
r0[53]=10'b1001001110;
r0[54]=10'b0001011110;
r0[55]=10'b1110001001;
r0[56]=10'b1110110001;
r0[57]=10'b1101111110;
r0[58]=10'b0111111000;
r0[59]=10'b1010001111;
r0[60]=10'b1100110100;
r0[61]=10'b0011010010;
r0[62]=10'b1101010100;
r0[63]=10'b1001110110;
//
r1[ 0]=10'b0100110000;
r1[ 1]=10'b0110000010;
r1[ 2]=10'b1110010001;
r1[ 3]=10'b0101110011;
r1[ 4]=10'b1011000110;
r1[ 5]=10'b1010101111;
r1[ 6]=10'b1110001000;
r1[ 7]=10'b0001010000;
r1[ 8]=10'b1011111100;
r1[ 9]=10'b0100010101;
r1[10]=10'b1100000100;
r1[11]=10'b0111011110;
r1[12]=10'b1001110011;
r1[13]=10'b1001101010;
r1[14]=10'b0001100101;
r1[15]=10'b0101101000;
r1[16]=10'b0111111011;
r1[17]=10'b1001110001;
r1[18]=10'b1101011001;
r1[19]=10'b0111011110;
r1[20]=10'b0011100101;
r1[21]=10'b1101000001;
r1[22]=10'b0110110001;
r1[23]=10'b0011000001;
r1[24]=10'b1111100001;
r1[25]=10'b0010011011;
r1[26]=10'b0110011110;
r1[27]=10'b0000111000;
r1[28]=10'b0000000101;
r1[29]=10'b0000100100;
r1[30]=10'b0110101101;
r1[31]=10'b1011010001;
r1[32]=10'b0001110111;
r1[33]=10'b0110100111;
r1[34]=10'b0111010101;
r1[35]=10'b1110110101;
r1[36]=10'b1011110110;
r1[37]=10'b1011011010;
r1[38]=10'b1100101010;
r1[39]=10'b1101101111;
r1[40]=10'b1110011111;
r1[41]=10'b1000100000;
r1[42]=10'b0110000101;
r1[43]=10'b0101111101;
r1[44]=10'b0011110111;
r1[45]=10'b1010001010;
r1[46]=10'b1101000011;
r1[47]=10'b1101101101;
r1[48]=10'b1011101001;
r1[49]=10'b0100001100;
r1[50]=10'b1001100010;
r1[51]=10'b1100110011;
r1[52]=10'b0011110101;
r1[53]=10'b0100110100;
r1[54]=10'b1110011000;
r1[55]=10'b1000111100;
r1[56]=10'b0100010000;
r1[57]=10'b0010011101;
r1[58]=10'b1100011010;
r1[59]=10'b0010011000;
r1[60]=10'b0001001000;
r1[61]=10'b0110001110;
r1[62]=10'b0110101101;
r1[63]=10'b1100011011; 
//

//
#5 ;
i=0;
end 
  // Update inputs on every positive edge of the clock
  always @(posedge clk_tb) begin
    if (i < 64) begin
      ao = r0[i];
      bo = r1[i];
      i = i + 1;
    end else begin
      #20; // Wait for some time before finishing the simulation
      $finish;
    end
  end


endmodule