module PRN_tb;
  reg clk_tb;
  reg [0:54] a, b;
  reg [0:4] c;
  wire [0:10229] p;
  wire [0:23] f, l;
reg  [0:54]r0[0:64];
reg [0:54]r1[0:64];
reg [0:5]c_1[0:64];
integer i;

  PRN P(.clk(clk_tb), .R0_in(a), .R1_in(b), .C_in(c), .P(p), .first(f), .last(l));

initial
begin
    clk_tb = 0;
end

always
begin
    #10;
    clk_tb = ~ clk_tb;
end


  initial begin
r0[0]=55'o0227743641272102303; 
r0[1]=55'o0603070242564637717;
r0[2]=55'o0746325144437416120;
r0[3]=55'o0023763714573206044;
r0[4]=55'o0155575663373106723;
r0[5]=55'o0022277536552741033;
r0[6]=55'o0137757627072411730;
r0[7]=55'o0413034001670700216;
r0[8]=55'o0501123675324707024;
r0[9]=55'o0013727517464264567;
r0[10]=55'o0663351450332761127;
r0[11]=55'o1450710073416110356;
r0[12]=55'o1716542347100366110;
r0[13]=55'o0743601273016301212;
r0[14]=55'o1454332372150500137;
r0[15]=55'o1473215015316613621;
r0[16]=55'o1255535602164437613;
r0[17]=55'o1164537254033266174;
r0[18]=55'o1500537251137244274;
r0[19]=55'o0766727150471256024;
r0[20]=55'o0457637114652202460;
r0[21]=55'o0436500136253056124;
r0[22]=55'o1666265767713037215;
r0[23]=55'o1465272157164065443;
r0[24]=55'o0607440357166466472;
r0[25]=55'o1670202421463640077;
r0[26]=55'o1312661744614412524;
r0[27]=55'o1413034001672741216;
r0[28]=55'o1113765722434040551;
r0[29]=55'o0621573414133237134;
r0[30]=55'o0526104310250410535;
r0[31]=55'o0426454733176070600;
r0[32]=55'o1440644676733136472;
r0[33]=55'o0557275325702027456;
r0[34]=55'o0657637150553356442;
r0[35]=55'o1403560400557766512;
r0[36]=55'o1531165662277124403;
r0[37]=55'o1403072012721162611;
r0[38]=55'o0541210077534050730;
r0[39]=55'o1660256422576622574;
r0[40]=55'o0646767375467672136;
r0[41]=55'o1563301635027210017;
r0[42]=55'o1403462012723163611;
r0[43]=55'o0767233376550711053;
r0[44]=55'o1260555130762307205;
r0[45]=55'o0531075060147161624;
r0[46]=55'o0112673710551347402;
r0[47]=55'o1314750013607403146;
r0[48]=55'o0471706447643213002;
r0[49]=55'o0770352206645261362;
r0[50]=55'o0255127616022236737;
r0[51]=55'o1035616240477274125;
r0[52]=55'o0251115713566666576;
r0[53]=55'o0752241454312660541;
r0[54]=55'o0461250256520434602;
r0[55]=55'o1116341217327713444;
r0[56]=55'o0765232132271554573;
r0[57]=55'o0774370107303671123;
r0[58]=55'o1407140711055577677;
r0[59]=55'o1753355476331367516;
r0[60]=55'o0101630163132222775;
r0[61]=55'o0730471404057577456;
r0[62]=55'o1336743247162047542;
r0[63]=55'o0020666576373544533;
//
r1[0]=55'o1667217344450257245 ;
r1[1]=55'o0300642746017221737 ;
r1[2]=55'o0474006332201753645 ;
r1[3]=55'o0613606702460402137 ;
r1[4]=55'o1465531713404064713 ;
r1[5]=55'o1063646422557130427 ;
r1[6]=55'o1066060465055002004 ;
r1[7]=55'o0225574416605070652 ;
r1[8]=55'o1733560674073230405 ;
r1[9]=55'o1116277147142260461 ;
r1[10]=55'o0663351450332761127 ;
r1[11]=55'o1110300535412261305 ;
r1[12]=55'o1046105227571557243 ;
r1[13]=55'o1020346561064461527 ;
r1[14]=55'o1270052747201123510 ;
r1[15]=55'o1041553307136735706 ;
r1[16]=55'o1002352163603013730 ;
r1[17]=55'o1362622514254366256 ;
r1[18]=55'o0556645716623157361 ;
r1[19]=55'o0020341533300021636 ;
r1[20]=55'o1470231623730254774 ;
r1[21]=55'o1437100574634755567 ;
r1[22]=55'o0215346037247347710 ;
r1[23]=55'o1074246275146357122 ;
r1[24]=55'o1655552356143710472 ;
r1[25]=55'o1067241424131022656 ;
r1[26]=55'o1611144345044137740 ;
r1[27]=55'o1235122601654653275 ;
r1[28]=55'o0663754302501454556 ;
r1[29]=55'o0330540311241344370 ;
r1[30]=55'o1763277034331577303 ;
r1[31]=55'o1325110610226320770 ;
r1[32]=55'o0632344657312671631 ;
r1[33]=55'o1432530060077160315 ;
r1[34]=55'o1272177170234542346 ;
r1[35]=55'o0043174152003062273 ;
r1[36]=55'o0633575650312403065 ;
r1[37]=55'o0305021033755066410 ;
r1[38]=55'o0137373436464572225 ;
r1[39]=55'o0014331642301151614 ;
r1[40]=55'o0444423305436737401 ;
r1[41]=55'o0232343171540161113 ;
r1[42]=55'o0101411166154322757 ;
r1[43]=55'o0501120665453153342 ;
r1[44]=55'o1042475051720150775 ;
r1[45]=55'o1533531265037673325 ;
r1[46]=55'o0506620200211067675 ;
r1[47]=55'o1324133406103765602 ;
r1[48]=55'o0203136107415235456 ;
r1[49]=55'o1521524233172031026 ;
r1[50]=55'o0164213410044443204 ;
r1[51]=55'o1221110757557452411 ;
r1[52]=55'o0252317630101475044 ;
r1[53]=55'o0014540074363706135 ;
r1[54]=55'o0371711523526255275 ;
r1[55]=55'o0012400567546521471 ;
r1[56]=55'o0312622351062337705 ;
r1[57]=55'o0023647344743400250 ;
r1[58]=55'o0257310611765747211 ;
r1[59]=55'o1540176212407214706 ;
r1[60]=55'o1412637164262406706 ;
r1[61]=55'o0363125736302421243 ;
r1[62]=55'o0414175374460515677 ;
r1[63]=55'o0004500310276201661 ;

c_1[0]=5'b01000 ;
c_1[1]=5'b00000 ;
c_1[2]=5'b01000 ;
c_1[3]=5'b00000 ;
c_1[4]=5'b01000 ;
c_1[5]=5'b01000 ;
c_1[6]=5'b00000 ;
c_1[7]=5'b01000 ;
c_1[8]=5'b00000 ;
c_1[9]=5'b00000 ;
c_1[10]=5'b00000 ;
c_1[11]=5'b01000 ;
c_1[12]=5'b01000 ;
c_1[13]=5'b00000 ;
c_1[14]=5'b00000 ;
c_1[15]=5'b00000 ;
c_1[16]=5'b01000 ;
c_1[17]=5'b01000 ;
c_1[18]=5'b01000 ;
c_1[19]=5'b01000 ;
c_1[20]=5'b00000 ;
c_1[21]=5'b01000 ;
c_1[22]=5'b01000 ;
c_1[23]=5'b00000 ;
c_1[24]=5'b01000 ;
c_1[25]=5'b00000 ;
c_1[26]=5'b01000 ;
c_1[27]=5'b00000 ;
c_1[28]=5'b00000 ;
c_1[29]=5'b00000 ;
c_1[30]=5'b00000 ;
c_1[31]=5'b01000 ;
c_1[32]=5'b01000 ;
c_1[33]=5'b00000 ;
c_1[34]=5'b01000 ;
c_1[35]=5'b01000 ;
c_1[36]=5'b00110 ;
c_1[37]=5'b00000 ;
c_1[38]=5'b01010 ;
c_1[39]=5'b00110 ;
c_1[40]=5'b00101 ;
c_1[41]=5'b10001 ;
c_1[42]=5'b00110 ;
c_1[43]=5'b00000 ;
c_1[44]=5'b10001 ;
c_1[45]=5'b00000 ;
c_1[46]=5'b00110 ;
c_1[47]=5'b00101 ;
c_1[48]=5'b00110 ;
c_1[49]=5'b10010 ;
c_1[50]=5'b10001 ;
c_1[51]=5'b00011 ;
c_1[52]=5'b01000 ;
c_1[53]=5'b00000 ;
c_1[54]=5'b00000 ;
c_1[55]=5'b00101 ;
c_1[56]=5'b10001 ;
c_1[57]=5'b00000 ;
c_1[58]=5'b01000 ;
c_1[59]=5'b00000 ;
c_1[60]=5'b00000 ;
c_1[61]=5'b10001 ;
c_1[62]=5'b00000 ;
c_1[63]=5'b01000 ;

#10 ;
i=0;
end 
  // Update inputs on every positive edge of the clock
  always @(posedge clk_tb) begin
    if (i < 64) begin
      a = r0[i];
      b = r1[i];
      c = c_1[i];
      i = i + 1;
    end else begin
      #20; // Wait for some time before finishing the simulation
      $finish;
    end
  end


endmodule







