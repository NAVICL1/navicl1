module PRN_tb2;
  reg clk_tb;
  reg [0:54] a2, b2;
  reg [0:4] c2;
  wire [0:10229] p2;
  wire [0:23] f2, l2;
reg  [0:54]r0[0:64];
reg [0:54]r1[0:64];
reg [0:54]c_1[0:64];
integer i;

  PRN P(.clk(clk_tb), .R0_in(a2), .R1_in(b2), .C_in(c2), .P(p2), .first(f2), .last(l2));

initial
begin
    clk_tb = 0;
end

always
begin
    #10;
    clk_tb = ~ clk_tb;
end


  initial begin
r0[0 ]=55'o0061727026503255544;
r0[1 ]=55'o1660130752435362260;
r0[2 ]=55'o0676457016477551225;
r0[3 ]=55'o1763467705267605701;
r0[4 ]=55'o1614265052776007236;
r0[5 ]=55'o1446113457553463523;
r0[6 ]=55'o1467417471470124574;
r0[7 ]=55'o0022513456555401603;
r0[8 ]=55'o0004420115402210365;
r0[9 ]=55'o0072276243316574510;
r0[10]=55'o1632356715721616750;
r0[11]=55'o1670164755420300763;
r0[12]=55'o1752127524253360255;
r0[13]=55'o0262220014044243135;
r0[14]=55'o1476157654546440020;
r0[15]=55'o1567545246612304745;
r0[16]=55'o0341667641424721673;
r0[17]=55'o0627234635353763045;
r0[18]=55'o0422600144741165152;
r0[19]=55'o1661124176724621030;
r0[20]=55'o1225124173720602330;
r0[21]=55'o1271773065617322065;
r0[22]=55'o0611751161355750124;
r0[23]=55'o0121046615341766266;
r0[24]=55'o0337423707274604122;
r0[25]=55'o0246610305446052270;
r0[26]=55'o0427326063324033344;
r0[27]=55'o1127467544162733403;
r0[28]=55'o0772425336125565156;
r0[29]=55'o1652465113031101044;
r0[30]=55'o1737622607214524550;
r0[31]=55'o1621315362240732407;
r0[32]=55'o0171733204500613155;
r0[33]=55'o1462031354327077565;
r0[34]=55'o1141265411761074755;
r0[35]=55'o0665106277260231251;
r0[36]=55'o0573123144343776027;
r0[37]=55'o0222101406610314705;
r0[38]=55'o0140673225434336401;
r0[39]=55'o0624233245727625631;
r0[40]=55'o0224022145647544263;
r0[41]=55'o0222501602610354705;
r0[42]=55'o1370337660412244327;
r0[43]=55'o0563567347256715524;
r0[44]=55'o1407636661116077143;
r0[45]=55'o1137431557133151004;
r0[46]=55'o1113003456475500265;
r0[47]=55'o1746553632646152413;
r0[48]=55'o1465416631251321074;
r0[49]=55'o0130516430377202712;
r0[50]=55'o0762173527246302776;
r0[51]=55'o1606732407336425136;
r0[52]=55'o1131112010066741562;
r0[53]=55'o1107467740060732403;
r0[54]=55'o0755500241327076744;
r0[55]=55'o1443037764170374631;
r0[56]=55'o0243224434357700345;
r0[57]=55'o0445504023027564357;
r0[58]=55'o1211152271373271472;
r0[59]=55'o0256644102553071753;
r0[60]=55'o0733312314424771412;
r0[61]=55'o1636376400221406415;
r0[62]=55'o0574114621235461516;
r0[63]=55'o1710717574016037362; 
//
r1[ 0]=55'o0377627103341647600;
r1[ 1]=55'o0047555332635133703;
r1[ 2]=55'o0570574070736102152;
r1[ 3]=55'o0511013576745450615;
r1[ 4]=55'o1216243446624447775;
r1[ 5]=55'o0176452272675511054;
r1[ 6]=55'o0151055342317137706;
r1[ 7]=55'o1127720116046071664;
r1[ 8]=55'o0514407436155575524;
r1[ 9]=55'o0253070462740453542;
r1[10]=55'o0573371306324706336;
r1[11]=55'o1315135317732077306;
r1[12]=55'o1170303027726635012;
r1[13]=55'o1637171270537414673;
r1[14]=55'o0342370520251732111;
r1[15]=55'o0142423551056551362;
r1[16]=55'o0641261355426453710;
r1[17]=55'o0237176034757345266;
r1[18]=55'o1205663360515365064;
r1[19]=55'o0725000004121104102;
r1[20]=55'o0337367500320303262;
r1[21]=55'o1303374445022536530;
r1[22]=55'o1033071464007363115;
r1[23]=55'o0753124124237073577;
r1[24]=55'o0133522075443754772;
r1[25]=55'o1244212514312345145;
r1[26]=55'o1066056211234322164;
r1[27]=55'o0073115240113351010;
r1[28]=55'o1102260031574577224;
r1[29]=55'o1166703527236520553;
r1[30]=55'o0056062273631723177;
r1[31]=55'o0141517013160576212;
r1[32]=55'o1644007677312431616;
r1[33]=55'o0201757033615262622;
r1[34]=55'o0357610362675720200;
r1[35]=55'o1637504174727237065;
r1[36]=55'o1510345507743707753;
r1[37]=55'o0540160763721100120;
r1[38]=55'o0406415410457500342;
r1[39]=55'o0707515543554212732;
r1[40]=55'o0140216674314371011;
r1[41]=55'o0445414471314273300;
r1[42]=55'o0120121661750263177;
r1[43]=55'o0477301251340044262;
r1[44]=55'o1157040657040363676;
r1[45]=55'o1222265021477405004;
r1[46]=55'o0314661556545362364;
r1[47]=55'o0177320240371640542;
r1[48]=55'o0735517310345570340;
r1[49]=55'o1367565551220511432;
r1[50]=55'o1274167141162675644;
r1[51]=55'o1543641015130470077;
r1[52]=55'o0640733734534576460;
r1[53]=55'o0216312531021205434;
r1[54]=55'o0050232164401566177;
r1[55]=55'o0702636370401726111;
r1[56]=55'o1733537351460015703;
r1[57]=55'o1523265651140460620;
r1[58]=55'o0607703231502460135;
r1[59]=55'o1757246242710445777;
r1[60]=55'o0464412467237572274;
r1[61]=55'o1050617751566552643;
r1[62]=55'o1041606123021052264;
r1[63]=55'o1335441345250455042;
//
c_1[ 0]=5'b10100;
c_1[ 1]=5'b10100;
c_1[ 2]=5'b00110;
c_1[ 3]=5'b10100;
c_1[ 4]=5'b10100;
c_1[ 5]=5'b00110;
c_1[ 6]=5'b10100;
c_1[ 7]=5'b00110;
c_1[ 8]=5'b00110;
c_1[ 9]=5'b00110;
c_1[10]=5'b10100;
c_1[11]=5'b00110;
c_1[12]=5'b10100;
c_1[13]=5'b00110;
c_1[14]=5'b00110;
c_1[15]=5'b10100;
c_1[16]=5'b00110;
c_1[17]=5'b00110;
c_1[18]=5'b00110;
c_1[19]=5'b00110;
c_1[20]=5'b10100;
c_1[21]=5'b10100;
c_1[22]=5'b10100;
c_1[23]=5'b00110;
c_1[24]=5'b10100;
c_1[25]=5'b00110;
c_1[26]=5'b00110;
c_1[27]=5'b00110;
c_1[28]=5'b00110;
c_1[29]=5'b10100;
c_1[30]=5'b10100;
c_1[31]=5'b00110;
c_1[32]=5'b10100;
c_1[33]=5'b00110;
c_1[34]=5'b00110;
c_1[35]=5'b00110;
c_1[36]=5'b10100;
c_1[37]=5'b10100;
c_1[38]=5'b01100;
c_1[39]=5'b00110;
c_1[40]=5'b00011;
c_1[41]=5'b01100;
c_1[42]=5'b10100;
c_1[43]=5'b00110;
c_1[44]=5'b10100;
c_1[45]=5'b10100;
c_1[46]=5'b00110;
c_1[47]=5'b00110;
c_1[48]=5'b00110;
c_1[49]=5'b10100;
c_1[50]=5'b10100;
c_1[51]=5'b10100;
c_1[52]=5'b00110;
c_1[53]=5'b10100;
c_1[54]=5'b00110;
c_1[55]=5'b10100;
c_1[56]=5'b00110;
c_1[57]=5'b00110;
c_1[58]=5'b10100;
c_1[59]=5'b10010;
c_1[60]=5'b10001;
c_1[61]=5'b11000;
c_1[62]=5'b00110;
c_1[63]=5'b10100;
//
#10 ;
i=0;
end 
  // Update inputs on every positive edge of the clock
  always @(posedge clk_tb) begin
    if (i < 64) begin
      a2 = r0[i];
      b2 = r1[i];
      c2 = c_1[i];
      i = i + 1;
    end else begin
      #20; // Wait for some time before finishing the simulation
      $finish;
    end
  end


endmodule
